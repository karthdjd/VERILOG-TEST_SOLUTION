module and_g_lev(input a,input b,output c);
  and(c,a,b);
endmodule
