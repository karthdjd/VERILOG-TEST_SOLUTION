module tristate_buff(input d,en,output y);
buf(y,d,en);
endmodule
